
`define USE_SRAM
`define SRAM_HEX_SIZE 7862
`define CRM_HEX_SIZE 0
`define DRAM_HEX_SIZE 0
`define HEX_SIZE 7862